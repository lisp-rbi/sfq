@SSR0F	CGTGCC	GHZ!Rj
@SSR1F	ATGCGT	GFHGGU