>My headerF
ATGCGTAGCGTAGCGATCGCTTCGTCGCTGTCGCTCGC
>mY headF
AAAAAAAAAAAAAAAATTTTTTTTTTTTTTTTGGGGGGGGG
