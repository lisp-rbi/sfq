>My header
ATGCGTAGCGTAGCGATCGCTTCGTCGCTGTCGCTCGC
>mY head
AAAAAAAAAAAAAAAATTTTTTTTTTTTTTTTGGGGGGGGG