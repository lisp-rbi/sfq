GHZ!Rj	@SSR0F	CGTGCC
GFHGGU	@SSR1F	ATGCGT